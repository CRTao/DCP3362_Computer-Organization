//Subject:     CO project 2 - Sign extend
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      
//----------------------------------------------
//Date:        
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------

module Sign_Extend(
    data_i,
    data_o
    );
               
//I/O ports
input   [16-1:0] data_i;
output  [32-1:0] data_o;

//Internal Signals
reg     [32-1:0] data_o;

//Sign extended

always @(*)begin
    data_o[32-1:16] = (data_i[16-1] == 1'b1) ? 16'b1111_1111_1111_1111:16'b0;
    data_o[16-1: 0] = data_i[16-1:0];
end         
		  
endmodule      
     